module Hex2SevenSeg(

	//////////// SEG7 //////////
	output	reg	     [7:0]		HEX,

	
	input 		     [3:0]		num
	
);

	always begin

	case (num)
		
		4'b0000: HEX[7:0] = 8'b11000000;
		4'b0001: HEX[7:0] = 8'b11111001;
		4'b0010: HEX[7:0] = 8'b10100100;
		4'b0011: HEX[7:0] = 8'b10110000;
		4'b0100: HEX[7:0] = 8'b10011001;
		4'b0101: HEX[7:0] = 8'b10010010;
		4'b0110: HEX[7:0] = 8'b10000010;
		4'b0111: HEX[7:0] = 8'b11111000;
		4'b1000: HEX[7:0] = 8'b10000000;
		4'b1001: HEX[7:0] = 8'b10010000;
		4'b1010: HEX[7:0] = 8'b10001000;
		4'b1011: HEX[7:0] = 8'b10000011;
		4'b1100: HEX[7:0] = 8'b11000110;
		4'b1101: HEX[7:0] = 8'b10100001;
		4'b1110: HEX[7:0] = 8'b10000110;
		4'b1111: HEX[7:0] = 8'b10001110;
      
      default : HEX[7:0] = 8'b11111111; // Default all segments off
		
		
	endcase







	end





endmodule